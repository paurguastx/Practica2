LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY GXOR IS
PORT( A, B: IN STD_LOGIC;
      X: OUT STD_LOGIC);
END GXOR;

ARCHITECTURE BEH OF GXOR IS
BEGIN
  X <= A XOR B;
END BEH;
